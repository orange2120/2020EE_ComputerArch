module HW4(clk,
            rst_n,
            // for mem_I
            mem_addr_I,
            mem_rdata_I,
			// for result output
			ctrl_signal,
			immediate,
			);

    input         clk, rst_n        ;
    output [31:2] mem_addr_I        ;
    input  [31:0] mem_rdata_I       ;
	output [11:0] ctrl_signal  ;
	output [31:0] immediate;
    
	// wire/reg 
	
	
	
	// Connect to your HW3 module


endmodule